module Memory(
  input        clock,
  input  [4:0] io_rdAddr,
  output [7:0] io_rdData,
  input        io_wrEna,
  input  [7:0] io_wrData,
  input  [4:0] io_wrAddr
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
  reg [7:0] mem [0:31]; // @[Memory.scala 16:16]
  wire [7:0] mem_io_rdData_MPORT_data; // @[Memory.scala 16:16]
  wire [4:0] mem_io_rdData_MPORT_addr; // @[Memory.scala 16:16]
  wire [7:0] mem_MPORT_data; // @[Memory.scala 16:16]
  wire [4:0] mem_MPORT_addr; // @[Memory.scala 16:16]
  wire  mem_MPORT_mask; // @[Memory.scala 16:16]
  wire  mem_MPORT_en; // @[Memory.scala 16:16]
  assign mem_io_rdData_MPORT_addr = io_rdAddr;
  assign mem_io_rdData_MPORT_data = mem[mem_io_rdData_MPORT_addr]; // @[Memory.scala 16:16]
  assign mem_MPORT_data = io_wrData;
  assign mem_MPORT_addr = io_wrAddr;
  assign mem_MPORT_mask = 1'h1;
  assign mem_MPORT_en = io_wrEna;
  assign io_rdData = mem_io_rdData_MPORT_data; // @[Memory.scala 25:13]
  always @(posedge clock) begin
    if(mem_MPORT_en & mem_MPORT_mask) begin
      mem[mem_MPORT_addr] <= mem_MPORT_data; // @[Memory.scala 16:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    mem[initvar] = _RAND_0[7:0];
`endif // RANDOMIZE_MEM_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module LiveValueTable(
  input        clock,
  input        reset,
  input  [4:0] io_wrAddr_0,
  input  [4:0] io_wrAddr_1,
  input  [4:0] io_wrAddr_2,
  input        io_wrEna_0,
  input        io_wrEna_1,
  input        io_wrEna_2,
  input  [4:0] io_rdAddr_0,
  input  [4:0] io_rdAddr_1,
  input  [4:0] io_rdAddr_2,
  output [1:0] io_rdIdx_0,
  output [1:0] io_rdIdx_1,
  output [1:0] io_rdIdx_2
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] lvtReg_0; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_1; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_2; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_3; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_4; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_5; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_6; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_7; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_8; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_9; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_10; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_11; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_12; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_13; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_14; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_15; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_16; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_17; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_18; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_19; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_20; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_21; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_22; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_23; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_24; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_25; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_26; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_27; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_28; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_29; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_30; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_31; // @[LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_0 = 5'h0 == io_wrAddr_0 ? 2'h0 : lvtReg_0; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1 = 5'h1 == io_wrAddr_0 ? 2'h0 : lvtReg_1; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_2 = 5'h2 == io_wrAddr_0 ? 2'h0 : lvtReg_2; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_3 = 5'h3 == io_wrAddr_0 ? 2'h0 : lvtReg_3; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_4 = 5'h4 == io_wrAddr_0 ? 2'h0 : lvtReg_4; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_5 = 5'h5 == io_wrAddr_0 ? 2'h0 : lvtReg_5; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_6 = 5'h6 == io_wrAddr_0 ? 2'h0 : lvtReg_6; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_7 = 5'h7 == io_wrAddr_0 ? 2'h0 : lvtReg_7; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_8 = 5'h8 == io_wrAddr_0 ? 2'h0 : lvtReg_8; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_9 = 5'h9 == io_wrAddr_0 ? 2'h0 : lvtReg_9; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_10 = 5'ha == io_wrAddr_0 ? 2'h0 : lvtReg_10; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_11 = 5'hb == io_wrAddr_0 ? 2'h0 : lvtReg_11; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_12 = 5'hc == io_wrAddr_0 ? 2'h0 : lvtReg_12; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_13 = 5'hd == io_wrAddr_0 ? 2'h0 : lvtReg_13; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_14 = 5'he == io_wrAddr_0 ? 2'h0 : lvtReg_14; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_15 = 5'hf == io_wrAddr_0 ? 2'h0 : lvtReg_15; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_16 = 5'h10 == io_wrAddr_0 ? 2'h0 : lvtReg_16; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_17 = 5'h11 == io_wrAddr_0 ? 2'h0 : lvtReg_17; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_18 = 5'h12 == io_wrAddr_0 ? 2'h0 : lvtReg_18; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_19 = 5'h13 == io_wrAddr_0 ? 2'h0 : lvtReg_19; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_20 = 5'h14 == io_wrAddr_0 ? 2'h0 : lvtReg_20; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_21 = 5'h15 == io_wrAddr_0 ? 2'h0 : lvtReg_21; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_22 = 5'h16 == io_wrAddr_0 ? 2'h0 : lvtReg_22; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_23 = 5'h17 == io_wrAddr_0 ? 2'h0 : lvtReg_23; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_24 = 5'h18 == io_wrAddr_0 ? 2'h0 : lvtReg_24; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_25 = 5'h19 == io_wrAddr_0 ? 2'h0 : lvtReg_25; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_26 = 5'h1a == io_wrAddr_0 ? 2'h0 : lvtReg_26; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_27 = 5'h1b == io_wrAddr_0 ? 2'h0 : lvtReg_27; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_28 = 5'h1c == io_wrAddr_0 ? 2'h0 : lvtReg_28; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_29 = 5'h1d == io_wrAddr_0 ? 2'h0 : lvtReg_29; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_30 = 5'h1e == io_wrAddr_0 ? 2'h0 : lvtReg_30; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_31 = 5'h1f == io_wrAddr_0 ? 2'h0 : lvtReg_31; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_32 = io_wrEna_0 ? _GEN_0 : lvtReg_0; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_33 = io_wrEna_0 ? _GEN_1 : lvtReg_1; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_34 = io_wrEna_0 ? _GEN_2 : lvtReg_2; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_35 = io_wrEna_0 ? _GEN_3 : lvtReg_3; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_36 = io_wrEna_0 ? _GEN_4 : lvtReg_4; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_37 = io_wrEna_0 ? _GEN_5 : lvtReg_5; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_38 = io_wrEna_0 ? _GEN_6 : lvtReg_6; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_39 = io_wrEna_0 ? _GEN_7 : lvtReg_7; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_40 = io_wrEna_0 ? _GEN_8 : lvtReg_8; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_41 = io_wrEna_0 ? _GEN_9 : lvtReg_9; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_42 = io_wrEna_0 ? _GEN_10 : lvtReg_10; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_43 = io_wrEna_0 ? _GEN_11 : lvtReg_11; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_44 = io_wrEna_0 ? _GEN_12 : lvtReg_12; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_45 = io_wrEna_0 ? _GEN_13 : lvtReg_13; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_46 = io_wrEna_0 ? _GEN_14 : lvtReg_14; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_47 = io_wrEna_0 ? _GEN_15 : lvtReg_15; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_48 = io_wrEna_0 ? _GEN_16 : lvtReg_16; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_49 = io_wrEna_0 ? _GEN_17 : lvtReg_17; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_50 = io_wrEna_0 ? _GEN_18 : lvtReg_18; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_51 = io_wrEna_0 ? _GEN_19 : lvtReg_19; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_52 = io_wrEna_0 ? _GEN_20 : lvtReg_20; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_53 = io_wrEna_0 ? _GEN_21 : lvtReg_21; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_54 = io_wrEna_0 ? _GEN_22 : lvtReg_22; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_55 = io_wrEna_0 ? _GEN_23 : lvtReg_23; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_56 = io_wrEna_0 ? _GEN_24 : lvtReg_24; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_57 = io_wrEna_0 ? _GEN_25 : lvtReg_25; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_58 = io_wrEna_0 ? _GEN_26 : lvtReg_26; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_59 = io_wrEna_0 ? _GEN_27 : lvtReg_27; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_60 = io_wrEna_0 ? _GEN_28 : lvtReg_28; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_61 = io_wrEna_0 ? _GEN_29 : lvtReg_29; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_62 = io_wrEna_0 ? _GEN_30 : lvtReg_30; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_63 = io_wrEna_0 ? _GEN_31 : lvtReg_31; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_64 = 5'h0 == io_wrAddr_1 ? 2'h1 : _GEN_32; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28]
  wire [1:0] _GEN_65 = 5'h1 == io_wrAddr_1 ? 2'h1 : _GEN_33; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28]
  wire [1:0] _GEN_66 = 5'h2 == io_wrAddr_1 ? 2'h1 : _GEN_34; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28]
  wire [1:0] _GEN_67 = 5'h3 == io_wrAddr_1 ? 2'h1 : _GEN_35; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28]
  wire [1:0] _GEN_68 = 5'h4 == io_wrAddr_1 ? 2'h1 : _GEN_36; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28]
  wire [1:0] _GEN_69 = 5'h5 == io_wrAddr_1 ? 2'h1 : _GEN_37; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28]
  wire [1:0] _GEN_70 = 5'h6 == io_wrAddr_1 ? 2'h1 : _GEN_38; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28]
  wire [1:0] _GEN_71 = 5'h7 == io_wrAddr_1 ? 2'h1 : _GEN_39; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28]
  wire [1:0] _GEN_72 = 5'h8 == io_wrAddr_1 ? 2'h1 : _GEN_40; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28]
  wire [1:0] _GEN_73 = 5'h9 == io_wrAddr_1 ? 2'h1 : _GEN_41; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28]
  wire [1:0] _GEN_74 = 5'ha == io_wrAddr_1 ? 2'h1 : _GEN_42; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28]
  wire [1:0] _GEN_75 = 5'hb == io_wrAddr_1 ? 2'h1 : _GEN_43; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28]
  wire [1:0] _GEN_76 = 5'hc == io_wrAddr_1 ? 2'h1 : _GEN_44; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28]
  wire [1:0] _GEN_77 = 5'hd == io_wrAddr_1 ? 2'h1 : _GEN_45; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28]
  wire [1:0] _GEN_78 = 5'he == io_wrAddr_1 ? 2'h1 : _GEN_46; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28]
  wire [1:0] _GEN_79 = 5'hf == io_wrAddr_1 ? 2'h1 : _GEN_47; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28]
  wire [1:0] _GEN_80 = 5'h10 == io_wrAddr_1 ? 2'h1 : _GEN_48; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28]
  wire [1:0] _GEN_81 = 5'h11 == io_wrAddr_1 ? 2'h1 : _GEN_49; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28]
  wire [1:0] _GEN_82 = 5'h12 == io_wrAddr_1 ? 2'h1 : _GEN_50; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28]
  wire [1:0] _GEN_83 = 5'h13 == io_wrAddr_1 ? 2'h1 : _GEN_51; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28]
  wire [1:0] _GEN_84 = 5'h14 == io_wrAddr_1 ? 2'h1 : _GEN_52; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28]
  wire [1:0] _GEN_85 = 5'h15 == io_wrAddr_1 ? 2'h1 : _GEN_53; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28]
  wire [1:0] _GEN_86 = 5'h16 == io_wrAddr_1 ? 2'h1 : _GEN_54; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28]
  wire [1:0] _GEN_87 = 5'h17 == io_wrAddr_1 ? 2'h1 : _GEN_55; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28]
  wire [1:0] _GEN_88 = 5'h18 == io_wrAddr_1 ? 2'h1 : _GEN_56; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28]
  wire [1:0] _GEN_89 = 5'h19 == io_wrAddr_1 ? 2'h1 : _GEN_57; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28]
  wire [1:0] _GEN_90 = 5'h1a == io_wrAddr_1 ? 2'h1 : _GEN_58; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28]
  wire [1:0] _GEN_91 = 5'h1b == io_wrAddr_1 ? 2'h1 : _GEN_59; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28]
  wire [1:0] _GEN_92 = 5'h1c == io_wrAddr_1 ? 2'h1 : _GEN_60; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28]
  wire [1:0] _GEN_93 = 5'h1d == io_wrAddr_1 ? 2'h1 : _GEN_61; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28]
  wire [1:0] _GEN_94 = 5'h1e == io_wrAddr_1 ? 2'h1 : _GEN_62; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28]
  wire [1:0] _GEN_95 = 5'h1f == io_wrAddr_1 ? 2'h1 : _GEN_63; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28]
  wire [1:0] _GEN_96 = io_wrEna_1 ? _GEN_64 : _GEN_32; // @[LVTMultiPortRams.scala 31:34]
  wire [1:0] _GEN_97 = io_wrEna_1 ? _GEN_65 : _GEN_33; // @[LVTMultiPortRams.scala 31:34]
  wire [1:0] _GEN_98 = io_wrEna_1 ? _GEN_66 : _GEN_34; // @[LVTMultiPortRams.scala 31:34]
  wire [1:0] _GEN_99 = io_wrEna_1 ? _GEN_67 : _GEN_35; // @[LVTMultiPortRams.scala 31:34]
  wire [1:0] _GEN_100 = io_wrEna_1 ? _GEN_68 : _GEN_36; // @[LVTMultiPortRams.scala 31:34]
  wire [1:0] _GEN_101 = io_wrEna_1 ? _GEN_69 : _GEN_37; // @[LVTMultiPortRams.scala 31:34]
  wire [1:0] _GEN_102 = io_wrEna_1 ? _GEN_70 : _GEN_38; // @[LVTMultiPortRams.scala 31:34]
  wire [1:0] _GEN_103 = io_wrEna_1 ? _GEN_71 : _GEN_39; // @[LVTMultiPortRams.scala 31:34]
  wire [1:0] _GEN_104 = io_wrEna_1 ? _GEN_72 : _GEN_40; // @[LVTMultiPortRams.scala 31:34]
  wire [1:0] _GEN_105 = io_wrEna_1 ? _GEN_73 : _GEN_41; // @[LVTMultiPortRams.scala 31:34]
  wire [1:0] _GEN_106 = io_wrEna_1 ? _GEN_74 : _GEN_42; // @[LVTMultiPortRams.scala 31:34]
  wire [1:0] _GEN_107 = io_wrEna_1 ? _GEN_75 : _GEN_43; // @[LVTMultiPortRams.scala 31:34]
  wire [1:0] _GEN_108 = io_wrEna_1 ? _GEN_76 : _GEN_44; // @[LVTMultiPortRams.scala 31:34]
  wire [1:0] _GEN_109 = io_wrEna_1 ? _GEN_77 : _GEN_45; // @[LVTMultiPortRams.scala 31:34]
  wire [1:0] _GEN_110 = io_wrEna_1 ? _GEN_78 : _GEN_46; // @[LVTMultiPortRams.scala 31:34]
  wire [1:0] _GEN_111 = io_wrEna_1 ? _GEN_79 : _GEN_47; // @[LVTMultiPortRams.scala 31:34]
  wire [1:0] _GEN_112 = io_wrEna_1 ? _GEN_80 : _GEN_48; // @[LVTMultiPortRams.scala 31:34]
  wire [1:0] _GEN_113 = io_wrEna_1 ? _GEN_81 : _GEN_49; // @[LVTMultiPortRams.scala 31:34]
  wire [1:0] _GEN_114 = io_wrEna_1 ? _GEN_82 : _GEN_50; // @[LVTMultiPortRams.scala 31:34]
  wire [1:0] _GEN_115 = io_wrEna_1 ? _GEN_83 : _GEN_51; // @[LVTMultiPortRams.scala 31:34]
  wire [1:0] _GEN_116 = io_wrEna_1 ? _GEN_84 : _GEN_52; // @[LVTMultiPortRams.scala 31:34]
  wire [1:0] _GEN_117 = io_wrEna_1 ? _GEN_85 : _GEN_53; // @[LVTMultiPortRams.scala 31:34]
  wire [1:0] _GEN_118 = io_wrEna_1 ? _GEN_86 : _GEN_54; // @[LVTMultiPortRams.scala 31:34]
  wire [1:0] _GEN_119 = io_wrEna_1 ? _GEN_87 : _GEN_55; // @[LVTMultiPortRams.scala 31:34]
  wire [1:0] _GEN_120 = io_wrEna_1 ? _GEN_88 : _GEN_56; // @[LVTMultiPortRams.scala 31:34]
  wire [1:0] _GEN_121 = io_wrEna_1 ? _GEN_89 : _GEN_57; // @[LVTMultiPortRams.scala 31:34]
  wire [1:0] _GEN_122 = io_wrEna_1 ? _GEN_90 : _GEN_58; // @[LVTMultiPortRams.scala 31:34]
  wire [1:0] _GEN_123 = io_wrEna_1 ? _GEN_91 : _GEN_59; // @[LVTMultiPortRams.scala 31:34]
  wire [1:0] _GEN_124 = io_wrEna_1 ? _GEN_92 : _GEN_60; // @[LVTMultiPortRams.scala 31:34]
  wire [1:0] _GEN_125 = io_wrEna_1 ? _GEN_93 : _GEN_61; // @[LVTMultiPortRams.scala 31:34]
  wire [1:0] _GEN_126 = io_wrEna_1 ? _GEN_94 : _GEN_62; // @[LVTMultiPortRams.scala 31:34]
  wire [1:0] _GEN_127 = io_wrEna_1 ? _GEN_95 : _GEN_63; // @[LVTMultiPortRams.scala 31:34]
  wire [1:0] _GEN_193 = 5'h1 == io_rdAddr_0 ? lvtReg_1 : lvtReg_0; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_194 = 5'h2 == io_rdAddr_0 ? lvtReg_2 : _GEN_193; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_195 = 5'h3 == io_rdAddr_0 ? lvtReg_3 : _GEN_194; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_196 = 5'h4 == io_rdAddr_0 ? lvtReg_4 : _GEN_195; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_197 = 5'h5 == io_rdAddr_0 ? lvtReg_5 : _GEN_196; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_198 = 5'h6 == io_rdAddr_0 ? lvtReg_6 : _GEN_197; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_199 = 5'h7 == io_rdAddr_0 ? lvtReg_7 : _GEN_198; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_200 = 5'h8 == io_rdAddr_0 ? lvtReg_8 : _GEN_199; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_201 = 5'h9 == io_rdAddr_0 ? lvtReg_9 : _GEN_200; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_202 = 5'ha == io_rdAddr_0 ? lvtReg_10 : _GEN_201; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_203 = 5'hb == io_rdAddr_0 ? lvtReg_11 : _GEN_202; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_204 = 5'hc == io_rdAddr_0 ? lvtReg_12 : _GEN_203; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_205 = 5'hd == io_rdAddr_0 ? lvtReg_13 : _GEN_204; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_206 = 5'he == io_rdAddr_0 ? lvtReg_14 : _GEN_205; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_207 = 5'hf == io_rdAddr_0 ? lvtReg_15 : _GEN_206; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_208 = 5'h10 == io_rdAddr_0 ? lvtReg_16 : _GEN_207; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_209 = 5'h11 == io_rdAddr_0 ? lvtReg_17 : _GEN_208; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_210 = 5'h12 == io_rdAddr_0 ? lvtReg_18 : _GEN_209; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_211 = 5'h13 == io_rdAddr_0 ? lvtReg_19 : _GEN_210; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_212 = 5'h14 == io_rdAddr_0 ? lvtReg_20 : _GEN_211; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_213 = 5'h15 == io_rdAddr_0 ? lvtReg_21 : _GEN_212; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_214 = 5'h16 == io_rdAddr_0 ? lvtReg_22 : _GEN_213; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_215 = 5'h17 == io_rdAddr_0 ? lvtReg_23 : _GEN_214; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_216 = 5'h18 == io_rdAddr_0 ? lvtReg_24 : _GEN_215; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_217 = 5'h19 == io_rdAddr_0 ? lvtReg_25 : _GEN_216; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_218 = 5'h1a == io_rdAddr_0 ? lvtReg_26 : _GEN_217; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_219 = 5'h1b == io_rdAddr_0 ? lvtReg_27 : _GEN_218; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_220 = 5'h1c == io_rdAddr_0 ? lvtReg_28 : _GEN_219; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_221 = 5'h1d == io_rdAddr_0 ? lvtReg_29 : _GEN_220; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_222 = 5'h1e == io_rdAddr_0 ? lvtReg_30 : _GEN_221; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_225 = 5'h1 == io_rdAddr_1 ? lvtReg_1 : lvtReg_0; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_226 = 5'h2 == io_rdAddr_1 ? lvtReg_2 : _GEN_225; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_227 = 5'h3 == io_rdAddr_1 ? lvtReg_3 : _GEN_226; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_228 = 5'h4 == io_rdAddr_1 ? lvtReg_4 : _GEN_227; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_229 = 5'h5 == io_rdAddr_1 ? lvtReg_5 : _GEN_228; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_230 = 5'h6 == io_rdAddr_1 ? lvtReg_6 : _GEN_229; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_231 = 5'h7 == io_rdAddr_1 ? lvtReg_7 : _GEN_230; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_232 = 5'h8 == io_rdAddr_1 ? lvtReg_8 : _GEN_231; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_233 = 5'h9 == io_rdAddr_1 ? lvtReg_9 : _GEN_232; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_234 = 5'ha == io_rdAddr_1 ? lvtReg_10 : _GEN_233; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_235 = 5'hb == io_rdAddr_1 ? lvtReg_11 : _GEN_234; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_236 = 5'hc == io_rdAddr_1 ? lvtReg_12 : _GEN_235; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_237 = 5'hd == io_rdAddr_1 ? lvtReg_13 : _GEN_236; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_238 = 5'he == io_rdAddr_1 ? lvtReg_14 : _GEN_237; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_239 = 5'hf == io_rdAddr_1 ? lvtReg_15 : _GEN_238; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_240 = 5'h10 == io_rdAddr_1 ? lvtReg_16 : _GEN_239; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_241 = 5'h11 == io_rdAddr_1 ? lvtReg_17 : _GEN_240; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_242 = 5'h12 == io_rdAddr_1 ? lvtReg_18 : _GEN_241; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_243 = 5'h13 == io_rdAddr_1 ? lvtReg_19 : _GEN_242; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_244 = 5'h14 == io_rdAddr_1 ? lvtReg_20 : _GEN_243; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_245 = 5'h15 == io_rdAddr_1 ? lvtReg_21 : _GEN_244; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_246 = 5'h16 == io_rdAddr_1 ? lvtReg_22 : _GEN_245; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_247 = 5'h17 == io_rdAddr_1 ? lvtReg_23 : _GEN_246; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_248 = 5'h18 == io_rdAddr_1 ? lvtReg_24 : _GEN_247; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_249 = 5'h19 == io_rdAddr_1 ? lvtReg_25 : _GEN_248; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_250 = 5'h1a == io_rdAddr_1 ? lvtReg_26 : _GEN_249; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_251 = 5'h1b == io_rdAddr_1 ? lvtReg_27 : _GEN_250; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_252 = 5'h1c == io_rdAddr_1 ? lvtReg_28 : _GEN_251; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_253 = 5'h1d == io_rdAddr_1 ? lvtReg_29 : _GEN_252; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_254 = 5'h1e == io_rdAddr_1 ? lvtReg_30 : _GEN_253; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_257 = 5'h1 == io_rdAddr_2 ? lvtReg_1 : lvtReg_0; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_258 = 5'h2 == io_rdAddr_2 ? lvtReg_2 : _GEN_257; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_259 = 5'h3 == io_rdAddr_2 ? lvtReg_3 : _GEN_258; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_260 = 5'h4 == io_rdAddr_2 ? lvtReg_4 : _GEN_259; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_261 = 5'h5 == io_rdAddr_2 ? lvtReg_5 : _GEN_260; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_262 = 5'h6 == io_rdAddr_2 ? lvtReg_6 : _GEN_261; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_263 = 5'h7 == io_rdAddr_2 ? lvtReg_7 : _GEN_262; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_264 = 5'h8 == io_rdAddr_2 ? lvtReg_8 : _GEN_263; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_265 = 5'h9 == io_rdAddr_2 ? lvtReg_9 : _GEN_264; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_266 = 5'ha == io_rdAddr_2 ? lvtReg_10 : _GEN_265; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_267 = 5'hb == io_rdAddr_2 ? lvtReg_11 : _GEN_266; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_268 = 5'hc == io_rdAddr_2 ? lvtReg_12 : _GEN_267; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_269 = 5'hd == io_rdAddr_2 ? lvtReg_13 : _GEN_268; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_270 = 5'he == io_rdAddr_2 ? lvtReg_14 : _GEN_269; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_271 = 5'hf == io_rdAddr_2 ? lvtReg_15 : _GEN_270; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_272 = 5'h10 == io_rdAddr_2 ? lvtReg_16 : _GEN_271; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_273 = 5'h11 == io_rdAddr_2 ? lvtReg_17 : _GEN_272; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_274 = 5'h12 == io_rdAddr_2 ? lvtReg_18 : _GEN_273; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_275 = 5'h13 == io_rdAddr_2 ? lvtReg_19 : _GEN_274; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_276 = 5'h14 == io_rdAddr_2 ? lvtReg_20 : _GEN_275; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_277 = 5'h15 == io_rdAddr_2 ? lvtReg_21 : _GEN_276; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_278 = 5'h16 == io_rdAddr_2 ? lvtReg_22 : _GEN_277; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_279 = 5'h17 == io_rdAddr_2 ? lvtReg_23 : _GEN_278; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_280 = 5'h18 == io_rdAddr_2 ? lvtReg_24 : _GEN_279; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_281 = 5'h19 == io_rdAddr_2 ? lvtReg_25 : _GEN_280; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_282 = 5'h1a == io_rdAddr_2 ? lvtReg_26 : _GEN_281; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_283 = 5'h1b == io_rdAddr_2 ? lvtReg_27 : _GEN_282; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_284 = 5'h1c == io_rdAddr_2 ? lvtReg_28 : _GEN_283; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_285 = 5'h1d == io_rdAddr_2 ? lvtReg_29 : _GEN_284; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_286 = 5'h1e == io_rdAddr_2 ? lvtReg_30 : _GEN_285; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  assign io_rdIdx_0 = 5'h1f == io_rdAddr_0 ? lvtReg_31 : _GEN_222; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  assign io_rdIdx_1 = 5'h1f == io_rdAddr_1 ? lvtReg_31 : _GEN_254; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  assign io_rdIdx_2 = 5'h1f == io_rdAddr_2 ? lvtReg_31 : _GEN_286; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  always @(posedge clock) begin
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_0 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_2) begin // @[LVTMultiPortRams.scala 31:34]
      if (5'h0 == io_wrAddr_2) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_0 <= 2'h2; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_0 <= _GEN_96;
      end
    end else begin
      lvtReg_0 <= _GEN_96;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_1 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_2) begin // @[LVTMultiPortRams.scala 31:34]
      if (5'h1 == io_wrAddr_2) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_1 <= 2'h2; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_1 <= _GEN_97;
      end
    end else begin
      lvtReg_1 <= _GEN_97;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_2 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_2) begin // @[LVTMultiPortRams.scala 31:34]
      if (5'h2 == io_wrAddr_2) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_2 <= 2'h2; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_2 <= _GEN_98;
      end
    end else begin
      lvtReg_2 <= _GEN_98;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_3 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_2) begin // @[LVTMultiPortRams.scala 31:34]
      if (5'h3 == io_wrAddr_2) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_3 <= 2'h2; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_3 <= _GEN_99;
      end
    end else begin
      lvtReg_3 <= _GEN_99;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_4 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_2) begin // @[LVTMultiPortRams.scala 31:34]
      if (5'h4 == io_wrAddr_2) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_4 <= 2'h2; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_4 <= _GEN_100;
      end
    end else begin
      lvtReg_4 <= _GEN_100;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_5 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_2) begin // @[LVTMultiPortRams.scala 31:34]
      if (5'h5 == io_wrAddr_2) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_5 <= 2'h2; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_5 <= _GEN_101;
      end
    end else begin
      lvtReg_5 <= _GEN_101;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_6 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_2) begin // @[LVTMultiPortRams.scala 31:34]
      if (5'h6 == io_wrAddr_2) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_6 <= 2'h2; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_6 <= _GEN_102;
      end
    end else begin
      lvtReg_6 <= _GEN_102;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_7 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_2) begin // @[LVTMultiPortRams.scala 31:34]
      if (5'h7 == io_wrAddr_2) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_7 <= 2'h2; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_7 <= _GEN_103;
      end
    end else begin
      lvtReg_7 <= _GEN_103;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_8 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_2) begin // @[LVTMultiPortRams.scala 31:34]
      if (5'h8 == io_wrAddr_2) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_8 <= 2'h2; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_8 <= _GEN_104;
      end
    end else begin
      lvtReg_8 <= _GEN_104;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_9 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_2) begin // @[LVTMultiPortRams.scala 31:34]
      if (5'h9 == io_wrAddr_2) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_9 <= 2'h2; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_9 <= _GEN_105;
      end
    end else begin
      lvtReg_9 <= _GEN_105;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_10 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_2) begin // @[LVTMultiPortRams.scala 31:34]
      if (5'ha == io_wrAddr_2) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_10 <= 2'h2; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_10 <= _GEN_106;
      end
    end else begin
      lvtReg_10 <= _GEN_106;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_11 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_2) begin // @[LVTMultiPortRams.scala 31:34]
      if (5'hb == io_wrAddr_2) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_11 <= 2'h2; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_11 <= _GEN_107;
      end
    end else begin
      lvtReg_11 <= _GEN_107;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_12 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_2) begin // @[LVTMultiPortRams.scala 31:34]
      if (5'hc == io_wrAddr_2) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_12 <= 2'h2; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_12 <= _GEN_108;
      end
    end else begin
      lvtReg_12 <= _GEN_108;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_13 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_2) begin // @[LVTMultiPortRams.scala 31:34]
      if (5'hd == io_wrAddr_2) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_13 <= 2'h2; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_13 <= _GEN_109;
      end
    end else begin
      lvtReg_13 <= _GEN_109;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_14 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_2) begin // @[LVTMultiPortRams.scala 31:34]
      if (5'he == io_wrAddr_2) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_14 <= 2'h2; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_14 <= _GEN_110;
      end
    end else begin
      lvtReg_14 <= _GEN_110;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_15 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_2) begin // @[LVTMultiPortRams.scala 31:34]
      if (5'hf == io_wrAddr_2) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_15 <= 2'h2; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_15 <= _GEN_111;
      end
    end else begin
      lvtReg_15 <= _GEN_111;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_16 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_2) begin // @[LVTMultiPortRams.scala 31:34]
      if (5'h10 == io_wrAddr_2) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_16 <= 2'h2; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_16 <= _GEN_112;
      end
    end else begin
      lvtReg_16 <= _GEN_112;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_17 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_2) begin // @[LVTMultiPortRams.scala 31:34]
      if (5'h11 == io_wrAddr_2) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_17 <= 2'h2; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_17 <= _GEN_113;
      end
    end else begin
      lvtReg_17 <= _GEN_113;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_18 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_2) begin // @[LVTMultiPortRams.scala 31:34]
      if (5'h12 == io_wrAddr_2) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_18 <= 2'h2; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_18 <= _GEN_114;
      end
    end else begin
      lvtReg_18 <= _GEN_114;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_19 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_2) begin // @[LVTMultiPortRams.scala 31:34]
      if (5'h13 == io_wrAddr_2) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_19 <= 2'h2; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_19 <= _GEN_115;
      end
    end else begin
      lvtReg_19 <= _GEN_115;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_20 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_2) begin // @[LVTMultiPortRams.scala 31:34]
      if (5'h14 == io_wrAddr_2) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_20 <= 2'h2; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_20 <= _GEN_116;
      end
    end else begin
      lvtReg_20 <= _GEN_116;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_21 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_2) begin // @[LVTMultiPortRams.scala 31:34]
      if (5'h15 == io_wrAddr_2) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_21 <= 2'h2; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_21 <= _GEN_117;
      end
    end else begin
      lvtReg_21 <= _GEN_117;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_22 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_2) begin // @[LVTMultiPortRams.scala 31:34]
      if (5'h16 == io_wrAddr_2) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_22 <= 2'h2; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_22 <= _GEN_118;
      end
    end else begin
      lvtReg_22 <= _GEN_118;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_23 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_2) begin // @[LVTMultiPortRams.scala 31:34]
      if (5'h17 == io_wrAddr_2) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_23 <= 2'h2; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_23 <= _GEN_119;
      end
    end else begin
      lvtReg_23 <= _GEN_119;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_24 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_2) begin // @[LVTMultiPortRams.scala 31:34]
      if (5'h18 == io_wrAddr_2) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_24 <= 2'h2; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_24 <= _GEN_120;
      end
    end else begin
      lvtReg_24 <= _GEN_120;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_25 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_2) begin // @[LVTMultiPortRams.scala 31:34]
      if (5'h19 == io_wrAddr_2) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_25 <= 2'h2; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_25 <= _GEN_121;
      end
    end else begin
      lvtReg_25 <= _GEN_121;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_26 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_2) begin // @[LVTMultiPortRams.scala 31:34]
      if (5'h1a == io_wrAddr_2) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_26 <= 2'h2; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_26 <= _GEN_122;
      end
    end else begin
      lvtReg_26 <= _GEN_122;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_27 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_2) begin // @[LVTMultiPortRams.scala 31:34]
      if (5'h1b == io_wrAddr_2) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_27 <= 2'h2; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_27 <= _GEN_123;
      end
    end else begin
      lvtReg_27 <= _GEN_123;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_28 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_2) begin // @[LVTMultiPortRams.scala 31:34]
      if (5'h1c == io_wrAddr_2) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_28 <= 2'h2; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_28 <= _GEN_124;
      end
    end else begin
      lvtReg_28 <= _GEN_124;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_29 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_2) begin // @[LVTMultiPortRams.scala 31:34]
      if (5'h1d == io_wrAddr_2) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_29 <= 2'h2; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_29 <= _GEN_125;
      end
    end else begin
      lvtReg_29 <= _GEN_125;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_30 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_2) begin // @[LVTMultiPortRams.scala 31:34]
      if (5'h1e == io_wrAddr_2) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_30 <= 2'h2; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_30 <= _GEN_126;
      end
    end else begin
      lvtReg_30 <= _GEN_126;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_31 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_2) begin // @[LVTMultiPortRams.scala 31:34]
      if (5'h1f == io_wrAddr_2) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_31 <= 2'h2; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_31 <= _GEN_127;
      end
    end else begin
      lvtReg_31 <= _GEN_127;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  lvtReg_0 = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  lvtReg_1 = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  lvtReg_2 = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  lvtReg_3 = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  lvtReg_4 = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  lvtReg_5 = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  lvtReg_6 = _RAND_6[1:0];
  _RAND_7 = {1{`RANDOM}};
  lvtReg_7 = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  lvtReg_8 = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  lvtReg_9 = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  lvtReg_10 = _RAND_10[1:0];
  _RAND_11 = {1{`RANDOM}};
  lvtReg_11 = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  lvtReg_12 = _RAND_12[1:0];
  _RAND_13 = {1{`RANDOM}};
  lvtReg_13 = _RAND_13[1:0];
  _RAND_14 = {1{`RANDOM}};
  lvtReg_14 = _RAND_14[1:0];
  _RAND_15 = {1{`RANDOM}};
  lvtReg_15 = _RAND_15[1:0];
  _RAND_16 = {1{`RANDOM}};
  lvtReg_16 = _RAND_16[1:0];
  _RAND_17 = {1{`RANDOM}};
  lvtReg_17 = _RAND_17[1:0];
  _RAND_18 = {1{`RANDOM}};
  lvtReg_18 = _RAND_18[1:0];
  _RAND_19 = {1{`RANDOM}};
  lvtReg_19 = _RAND_19[1:0];
  _RAND_20 = {1{`RANDOM}};
  lvtReg_20 = _RAND_20[1:0];
  _RAND_21 = {1{`RANDOM}};
  lvtReg_21 = _RAND_21[1:0];
  _RAND_22 = {1{`RANDOM}};
  lvtReg_22 = _RAND_22[1:0];
  _RAND_23 = {1{`RANDOM}};
  lvtReg_23 = _RAND_23[1:0];
  _RAND_24 = {1{`RANDOM}};
  lvtReg_24 = _RAND_24[1:0];
  _RAND_25 = {1{`RANDOM}};
  lvtReg_25 = _RAND_25[1:0];
  _RAND_26 = {1{`RANDOM}};
  lvtReg_26 = _RAND_26[1:0];
  _RAND_27 = {1{`RANDOM}};
  lvtReg_27 = _RAND_27[1:0];
  _RAND_28 = {1{`RANDOM}};
  lvtReg_28 = _RAND_28[1:0];
  _RAND_29 = {1{`RANDOM}};
  lvtReg_29 = _RAND_29[1:0];
  _RAND_30 = {1{`RANDOM}};
  lvtReg_30 = _RAND_30[1:0];
  _RAND_31 = {1{`RANDOM}};
  lvtReg_31 = _RAND_31[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module LVTMultiPortRams(
  input        clock,
  input        reset,
  input  [4:0] io_wrAddr_0,
  input  [4:0] io_wrAddr_1,
  input  [4:0] io_wrAddr_2,
  input  [7:0] io_wrData_0,
  input  [7:0] io_wrData_1,
  input  [7:0] io_wrData_2,
  input        io_wrEna_0,
  input        io_wrEna_1,
  input        io_wrEna_2,
  input  [4:0] io_rdAddr_0,
  input  [4:0] io_rdAddr_1,
  input  [4:0] io_rdAddr_2,
  output [7:0] io_rdData_0,
  output [7:0] io_rdData_1,
  output [7:0] io_rdData_2
);
  wire  Memory_clock; // @[LVTMultiPortRams.scala 52:44]
  wire [4:0] Memory_io_rdAddr; // @[LVTMultiPortRams.scala 52:44]
  wire [7:0] Memory_io_rdData; // @[LVTMultiPortRams.scala 52:44]
  wire  Memory_io_wrEna; // @[LVTMultiPortRams.scala 52:44]
  wire [7:0] Memory_io_wrData; // @[LVTMultiPortRams.scala 52:44]
  wire [4:0] Memory_io_wrAddr; // @[LVTMultiPortRams.scala 52:44]
  wire  Memory_1_clock; // @[LVTMultiPortRams.scala 52:44]
  wire [4:0] Memory_1_io_rdAddr; // @[LVTMultiPortRams.scala 52:44]
  wire [7:0] Memory_1_io_rdData; // @[LVTMultiPortRams.scala 52:44]
  wire  Memory_1_io_wrEna; // @[LVTMultiPortRams.scala 52:44]
  wire [7:0] Memory_1_io_wrData; // @[LVTMultiPortRams.scala 52:44]
  wire [4:0] Memory_1_io_wrAddr; // @[LVTMultiPortRams.scala 52:44]
  wire  Memory_2_clock; // @[LVTMultiPortRams.scala 52:44]
  wire [4:0] Memory_2_io_rdAddr; // @[LVTMultiPortRams.scala 52:44]
  wire [7:0] Memory_2_io_rdData; // @[LVTMultiPortRams.scala 52:44]
  wire  Memory_2_io_wrEna; // @[LVTMultiPortRams.scala 52:44]
  wire [7:0] Memory_2_io_wrData; // @[LVTMultiPortRams.scala 52:44]
  wire [4:0] Memory_2_io_wrAddr; // @[LVTMultiPortRams.scala 52:44]
  wire  Memory_3_clock; // @[LVTMultiPortRams.scala 52:44]
  wire [4:0] Memory_3_io_rdAddr; // @[LVTMultiPortRams.scala 52:44]
  wire [7:0] Memory_3_io_rdData; // @[LVTMultiPortRams.scala 52:44]
  wire  Memory_3_io_wrEna; // @[LVTMultiPortRams.scala 52:44]
  wire [7:0] Memory_3_io_wrData; // @[LVTMultiPortRams.scala 52:44]
  wire [4:0] Memory_3_io_wrAddr; // @[LVTMultiPortRams.scala 52:44]
  wire  Memory_4_clock; // @[LVTMultiPortRams.scala 52:44]
  wire [4:0] Memory_4_io_rdAddr; // @[LVTMultiPortRams.scala 52:44]
  wire [7:0] Memory_4_io_rdData; // @[LVTMultiPortRams.scala 52:44]
  wire  Memory_4_io_wrEna; // @[LVTMultiPortRams.scala 52:44]
  wire [7:0] Memory_4_io_wrData; // @[LVTMultiPortRams.scala 52:44]
  wire [4:0] Memory_4_io_wrAddr; // @[LVTMultiPortRams.scala 52:44]
  wire  Memory_5_clock; // @[LVTMultiPortRams.scala 52:44]
  wire [4:0] Memory_5_io_rdAddr; // @[LVTMultiPortRams.scala 52:44]
  wire [7:0] Memory_5_io_rdData; // @[LVTMultiPortRams.scala 52:44]
  wire  Memory_5_io_wrEna; // @[LVTMultiPortRams.scala 52:44]
  wire [7:0] Memory_5_io_wrData; // @[LVTMultiPortRams.scala 52:44]
  wire [4:0] Memory_5_io_wrAddr; // @[LVTMultiPortRams.scala 52:44]
  wire  Memory_6_clock; // @[LVTMultiPortRams.scala 52:44]
  wire [4:0] Memory_6_io_rdAddr; // @[LVTMultiPortRams.scala 52:44]
  wire [7:0] Memory_6_io_rdData; // @[LVTMultiPortRams.scala 52:44]
  wire  Memory_6_io_wrEna; // @[LVTMultiPortRams.scala 52:44]
  wire [7:0] Memory_6_io_wrData; // @[LVTMultiPortRams.scala 52:44]
  wire [4:0] Memory_6_io_wrAddr; // @[LVTMultiPortRams.scala 52:44]
  wire  Memory_7_clock; // @[LVTMultiPortRams.scala 52:44]
  wire [4:0] Memory_7_io_rdAddr; // @[LVTMultiPortRams.scala 52:44]
  wire [7:0] Memory_7_io_rdData; // @[LVTMultiPortRams.scala 52:44]
  wire  Memory_7_io_wrEna; // @[LVTMultiPortRams.scala 52:44]
  wire [7:0] Memory_7_io_wrData; // @[LVTMultiPortRams.scala 52:44]
  wire [4:0] Memory_7_io_wrAddr; // @[LVTMultiPortRams.scala 52:44]
  wire  Memory_8_clock; // @[LVTMultiPortRams.scala 52:44]
  wire [4:0] Memory_8_io_rdAddr; // @[LVTMultiPortRams.scala 52:44]
  wire [7:0] Memory_8_io_rdData; // @[LVTMultiPortRams.scala 52:44]
  wire  Memory_8_io_wrEna; // @[LVTMultiPortRams.scala 52:44]
  wire [7:0] Memory_8_io_wrData; // @[LVTMultiPortRams.scala 52:44]
  wire [4:0] Memory_8_io_wrAddr; // @[LVTMultiPortRams.scala 52:44]
  wire  lvt_clock; // @[LVTMultiPortRams.scala 53:19]
  wire  lvt_reset; // @[LVTMultiPortRams.scala 53:19]
  wire [4:0] lvt_io_wrAddr_0; // @[LVTMultiPortRams.scala 53:19]
  wire [4:0] lvt_io_wrAddr_1; // @[LVTMultiPortRams.scala 53:19]
  wire [4:0] lvt_io_wrAddr_2; // @[LVTMultiPortRams.scala 53:19]
  wire  lvt_io_wrEna_0; // @[LVTMultiPortRams.scala 53:19]
  wire  lvt_io_wrEna_1; // @[LVTMultiPortRams.scala 53:19]
  wire  lvt_io_wrEna_2; // @[LVTMultiPortRams.scala 53:19]
  wire [4:0] lvt_io_rdAddr_0; // @[LVTMultiPortRams.scala 53:19]
  wire [4:0] lvt_io_rdAddr_1; // @[LVTMultiPortRams.scala 53:19]
  wire [4:0] lvt_io_rdAddr_2; // @[LVTMultiPortRams.scala 53:19]
  wire [1:0] lvt_io_rdIdx_0; // @[LVTMultiPortRams.scala 53:19]
  wire [1:0] lvt_io_rdIdx_1; // @[LVTMultiPortRams.scala 53:19]
  wire [1:0] lvt_io_rdIdx_2; // @[LVTMultiPortRams.scala 53:19]
  wire [3:0] _io_rdData_0_T = lvt_io_rdIdx_0 * 2'h3; // @[LVTMultiPortRams.scala 72:30]
  wire [4:0] _io_rdData_0_T_1 = {{1'd0}, _io_rdData_0_T}; // @[LVTMultiPortRams.scala 72:36]
  wire [7:0] mems_0_rdData = Memory_io_rdData; // @[LVTMultiPortRams.scala 52:21 LVTMultiPortRams.scala 52:21]
  wire [7:0] mems_1_rdData = Memory_1_io_rdData; // @[LVTMultiPortRams.scala 52:21 LVTMultiPortRams.scala 52:21]
  wire [7:0] _GEN_6 = 4'h1 == _io_rdData_0_T_1[3:0] ? mems_1_rdData : mems_0_rdData; // @[LVTMultiPortRams.scala 72:18 LVTMultiPortRams.scala 72:18]
  wire [7:0] mems_2_rdData = Memory_2_io_rdData; // @[LVTMultiPortRams.scala 52:21 LVTMultiPortRams.scala 52:21]
  wire [7:0] _GEN_11 = 4'h2 == _io_rdData_0_T_1[3:0] ? mems_2_rdData : _GEN_6; // @[LVTMultiPortRams.scala 72:18 LVTMultiPortRams.scala 72:18]
  wire [7:0] mems_3_rdData = Memory_3_io_rdData; // @[LVTMultiPortRams.scala 52:21 LVTMultiPortRams.scala 52:21]
  wire [7:0] _GEN_16 = 4'h3 == _io_rdData_0_T_1[3:0] ? mems_3_rdData : _GEN_11; // @[LVTMultiPortRams.scala 72:18 LVTMultiPortRams.scala 72:18]
  wire [7:0] mems_4_rdData = Memory_4_io_rdData; // @[LVTMultiPortRams.scala 52:21 LVTMultiPortRams.scala 52:21]
  wire [7:0] _GEN_21 = 4'h4 == _io_rdData_0_T_1[3:0] ? mems_4_rdData : _GEN_16; // @[LVTMultiPortRams.scala 72:18 LVTMultiPortRams.scala 72:18]
  wire [7:0] mems_5_rdData = Memory_5_io_rdData; // @[LVTMultiPortRams.scala 52:21 LVTMultiPortRams.scala 52:21]
  wire [7:0] _GEN_26 = 4'h5 == _io_rdData_0_T_1[3:0] ? mems_5_rdData : _GEN_21; // @[LVTMultiPortRams.scala 72:18 LVTMultiPortRams.scala 72:18]
  wire [7:0] mems_6_rdData = Memory_6_io_rdData; // @[LVTMultiPortRams.scala 52:21 LVTMultiPortRams.scala 52:21]
  wire [7:0] _GEN_31 = 4'h6 == _io_rdData_0_T_1[3:0] ? mems_6_rdData : _GEN_26; // @[LVTMultiPortRams.scala 72:18 LVTMultiPortRams.scala 72:18]
  wire [7:0] mems_7_rdData = Memory_7_io_rdData; // @[LVTMultiPortRams.scala 52:21 LVTMultiPortRams.scala 52:21]
  wire [7:0] _GEN_36 = 4'h7 == _io_rdData_0_T_1[3:0] ? mems_7_rdData : _GEN_31; // @[LVTMultiPortRams.scala 72:18 LVTMultiPortRams.scala 72:18]
  wire [7:0] mems_8_rdData = Memory_8_io_rdData; // @[LVTMultiPortRams.scala 52:21 LVTMultiPortRams.scala 52:21]
  wire [3:0] _io_rdData_1_T = lvt_io_rdIdx_1 * 2'h3; // @[LVTMultiPortRams.scala 72:30]
  wire [3:0] _io_rdData_1_T_2 = _io_rdData_1_T + 4'h1; // @[LVTMultiPortRams.scala 72:36]
  wire [7:0] _GEN_51 = 4'h1 == _io_rdData_1_T_2 ? mems_1_rdData : mems_0_rdData; // @[LVTMultiPortRams.scala 72:18 LVTMultiPortRams.scala 72:18]
  wire [7:0] _GEN_56 = 4'h2 == _io_rdData_1_T_2 ? mems_2_rdData : _GEN_51; // @[LVTMultiPortRams.scala 72:18 LVTMultiPortRams.scala 72:18]
  wire [7:0] _GEN_61 = 4'h3 == _io_rdData_1_T_2 ? mems_3_rdData : _GEN_56; // @[LVTMultiPortRams.scala 72:18 LVTMultiPortRams.scala 72:18]
  wire [7:0] _GEN_66 = 4'h4 == _io_rdData_1_T_2 ? mems_4_rdData : _GEN_61; // @[LVTMultiPortRams.scala 72:18 LVTMultiPortRams.scala 72:18]
  wire [7:0] _GEN_71 = 4'h5 == _io_rdData_1_T_2 ? mems_5_rdData : _GEN_66; // @[LVTMultiPortRams.scala 72:18 LVTMultiPortRams.scala 72:18]
  wire [7:0] _GEN_76 = 4'h6 == _io_rdData_1_T_2 ? mems_6_rdData : _GEN_71; // @[LVTMultiPortRams.scala 72:18 LVTMultiPortRams.scala 72:18]
  wire [7:0] _GEN_81 = 4'h7 == _io_rdData_1_T_2 ? mems_7_rdData : _GEN_76; // @[LVTMultiPortRams.scala 72:18 LVTMultiPortRams.scala 72:18]
  wire [3:0] _io_rdData_2_T = lvt_io_rdIdx_2 * 2'h3; // @[LVTMultiPortRams.scala 72:30]
  wire [3:0] _io_rdData_2_T_2 = _io_rdData_2_T + 4'h2; // @[LVTMultiPortRams.scala 72:36]
  wire [7:0] _GEN_96 = 4'h1 == _io_rdData_2_T_2 ? mems_1_rdData : mems_0_rdData; // @[LVTMultiPortRams.scala 72:18 LVTMultiPortRams.scala 72:18]
  wire [7:0] _GEN_101 = 4'h2 == _io_rdData_2_T_2 ? mems_2_rdData : _GEN_96; // @[LVTMultiPortRams.scala 72:18 LVTMultiPortRams.scala 72:18]
  wire [7:0] _GEN_106 = 4'h3 == _io_rdData_2_T_2 ? mems_3_rdData : _GEN_101; // @[LVTMultiPortRams.scala 72:18 LVTMultiPortRams.scala 72:18]
  wire [7:0] _GEN_111 = 4'h4 == _io_rdData_2_T_2 ? mems_4_rdData : _GEN_106; // @[LVTMultiPortRams.scala 72:18 LVTMultiPortRams.scala 72:18]
  wire [7:0] _GEN_116 = 4'h5 == _io_rdData_2_T_2 ? mems_5_rdData : _GEN_111; // @[LVTMultiPortRams.scala 72:18 LVTMultiPortRams.scala 72:18]
  wire [7:0] _GEN_121 = 4'h6 == _io_rdData_2_T_2 ? mems_6_rdData : _GEN_116; // @[LVTMultiPortRams.scala 72:18 LVTMultiPortRams.scala 72:18]
  wire [7:0] _GEN_126 = 4'h7 == _io_rdData_2_T_2 ? mems_7_rdData : _GEN_121; // @[LVTMultiPortRams.scala 72:18 LVTMultiPortRams.scala 72:18]
  Memory Memory ( // @[LVTMultiPortRams.scala 52:44]
    .clock(Memory_clock),
    .io_rdAddr(Memory_io_rdAddr),
    .io_rdData(Memory_io_rdData),
    .io_wrEna(Memory_io_wrEna),
    .io_wrData(Memory_io_wrData),
    .io_wrAddr(Memory_io_wrAddr)
  );
  Memory Memory_1 ( // @[LVTMultiPortRams.scala 52:44]
    .clock(Memory_1_clock),
    .io_rdAddr(Memory_1_io_rdAddr),
    .io_rdData(Memory_1_io_rdData),
    .io_wrEna(Memory_1_io_wrEna),
    .io_wrData(Memory_1_io_wrData),
    .io_wrAddr(Memory_1_io_wrAddr)
  );
  Memory Memory_2 ( // @[LVTMultiPortRams.scala 52:44]
    .clock(Memory_2_clock),
    .io_rdAddr(Memory_2_io_rdAddr),
    .io_rdData(Memory_2_io_rdData),
    .io_wrEna(Memory_2_io_wrEna),
    .io_wrData(Memory_2_io_wrData),
    .io_wrAddr(Memory_2_io_wrAddr)
  );
  Memory Memory_3 ( // @[LVTMultiPortRams.scala 52:44]
    .clock(Memory_3_clock),
    .io_rdAddr(Memory_3_io_rdAddr),
    .io_rdData(Memory_3_io_rdData),
    .io_wrEna(Memory_3_io_wrEna),
    .io_wrData(Memory_3_io_wrData),
    .io_wrAddr(Memory_3_io_wrAddr)
  );
  Memory Memory_4 ( // @[LVTMultiPortRams.scala 52:44]
    .clock(Memory_4_clock),
    .io_rdAddr(Memory_4_io_rdAddr),
    .io_rdData(Memory_4_io_rdData),
    .io_wrEna(Memory_4_io_wrEna),
    .io_wrData(Memory_4_io_wrData),
    .io_wrAddr(Memory_4_io_wrAddr)
  );
  Memory Memory_5 ( // @[LVTMultiPortRams.scala 52:44]
    .clock(Memory_5_clock),
    .io_rdAddr(Memory_5_io_rdAddr),
    .io_rdData(Memory_5_io_rdData),
    .io_wrEna(Memory_5_io_wrEna),
    .io_wrData(Memory_5_io_wrData),
    .io_wrAddr(Memory_5_io_wrAddr)
  );
  Memory Memory_6 ( // @[LVTMultiPortRams.scala 52:44]
    .clock(Memory_6_clock),
    .io_rdAddr(Memory_6_io_rdAddr),
    .io_rdData(Memory_6_io_rdData),
    .io_wrEna(Memory_6_io_wrEna),
    .io_wrData(Memory_6_io_wrData),
    .io_wrAddr(Memory_6_io_wrAddr)
  );
  Memory Memory_7 ( // @[LVTMultiPortRams.scala 52:44]
    .clock(Memory_7_clock),
    .io_rdAddr(Memory_7_io_rdAddr),
    .io_rdData(Memory_7_io_rdData),
    .io_wrEna(Memory_7_io_wrEna),
    .io_wrData(Memory_7_io_wrData),
    .io_wrAddr(Memory_7_io_wrAddr)
  );
  Memory Memory_8 ( // @[LVTMultiPortRams.scala 52:44]
    .clock(Memory_8_clock),
    .io_rdAddr(Memory_8_io_rdAddr),
    .io_rdData(Memory_8_io_rdData),
    .io_wrEna(Memory_8_io_wrEna),
    .io_wrData(Memory_8_io_wrData),
    .io_wrAddr(Memory_8_io_wrAddr)
  );
  LiveValueTable lvt ( // @[LVTMultiPortRams.scala 53:19]
    .clock(lvt_clock),
    .reset(lvt_reset),
    .io_wrAddr_0(lvt_io_wrAddr_0),
    .io_wrAddr_1(lvt_io_wrAddr_1),
    .io_wrAddr_2(lvt_io_wrAddr_2),
    .io_wrEna_0(lvt_io_wrEna_0),
    .io_wrEna_1(lvt_io_wrEna_1),
    .io_wrEna_2(lvt_io_wrEna_2),
    .io_rdAddr_0(lvt_io_rdAddr_0),
    .io_rdAddr_1(lvt_io_rdAddr_1),
    .io_rdAddr_2(lvt_io_rdAddr_2),
    .io_rdIdx_0(lvt_io_rdIdx_0),
    .io_rdIdx_1(lvt_io_rdIdx_1),
    .io_rdIdx_2(lvt_io_rdIdx_2)
  );
  assign io_rdData_0 = 4'h8 == _io_rdData_0_T_1[3:0] ? mems_8_rdData : _GEN_36; // @[LVTMultiPortRams.scala 72:18 LVTMultiPortRams.scala 72:18]
  assign io_rdData_1 = 4'h8 == _io_rdData_1_T_2 ? mems_8_rdData : _GEN_81; // @[LVTMultiPortRams.scala 72:18 LVTMultiPortRams.scala 72:18]
  assign io_rdData_2 = 4'h8 == _io_rdData_2_T_2 ? mems_8_rdData : _GEN_126; // @[LVTMultiPortRams.scala 72:18 LVTMultiPortRams.scala 72:18]
  assign Memory_clock = clock;
  assign Memory_io_rdAddr = io_rdAddr_0; // @[LVTMultiPortRams.scala 52:21 LVTMultiPortRams.scala 60:30]
  assign Memory_io_wrEna = io_wrEna_0; // @[LVTMultiPortRams.scala 52:21 LVTMultiPortRams.scala 57:29]
  assign Memory_io_wrData = io_wrData_0; // @[LVTMultiPortRams.scala 52:21 LVTMultiPortRams.scala 59:30]
  assign Memory_io_wrAddr = io_wrAddr_0; // @[LVTMultiPortRams.scala 52:21 LVTMultiPortRams.scala 58:30]
  assign Memory_1_clock = clock;
  assign Memory_1_io_rdAddr = io_rdAddr_1; // @[LVTMultiPortRams.scala 52:21 LVTMultiPortRams.scala 60:30]
  assign Memory_1_io_wrEna = io_wrEna_0; // @[LVTMultiPortRams.scala 52:21 LVTMultiPortRams.scala 57:29]
  assign Memory_1_io_wrData = io_wrData_0; // @[LVTMultiPortRams.scala 52:21 LVTMultiPortRams.scala 59:30]
  assign Memory_1_io_wrAddr = io_wrAddr_0; // @[LVTMultiPortRams.scala 52:21 LVTMultiPortRams.scala 58:30]
  assign Memory_2_clock = clock;
  assign Memory_2_io_rdAddr = io_rdAddr_2; // @[LVTMultiPortRams.scala 52:21 LVTMultiPortRams.scala 60:30]
  assign Memory_2_io_wrEna = io_wrEna_0; // @[LVTMultiPortRams.scala 52:21 LVTMultiPortRams.scala 57:29]
  assign Memory_2_io_wrData = io_wrData_0; // @[LVTMultiPortRams.scala 52:21 LVTMultiPortRams.scala 59:30]
  assign Memory_2_io_wrAddr = io_wrAddr_0; // @[LVTMultiPortRams.scala 52:21 LVTMultiPortRams.scala 58:30]
  assign Memory_3_clock = clock;
  assign Memory_3_io_rdAddr = io_rdAddr_0; // @[LVTMultiPortRams.scala 52:21 LVTMultiPortRams.scala 60:30]
  assign Memory_3_io_wrEna = io_wrEna_1; // @[LVTMultiPortRams.scala 52:21 LVTMultiPortRams.scala 57:29]
  assign Memory_3_io_wrData = io_wrData_1; // @[LVTMultiPortRams.scala 52:21 LVTMultiPortRams.scala 59:30]
  assign Memory_3_io_wrAddr = io_wrAddr_1; // @[LVTMultiPortRams.scala 52:21 LVTMultiPortRams.scala 58:30]
  assign Memory_4_clock = clock;
  assign Memory_4_io_rdAddr = io_rdAddr_1; // @[LVTMultiPortRams.scala 52:21 LVTMultiPortRams.scala 60:30]
  assign Memory_4_io_wrEna = io_wrEna_1; // @[LVTMultiPortRams.scala 52:21 LVTMultiPortRams.scala 57:29]
  assign Memory_4_io_wrData = io_wrData_1; // @[LVTMultiPortRams.scala 52:21 LVTMultiPortRams.scala 59:30]
  assign Memory_4_io_wrAddr = io_wrAddr_1; // @[LVTMultiPortRams.scala 52:21 LVTMultiPortRams.scala 58:30]
  assign Memory_5_clock = clock;
  assign Memory_5_io_rdAddr = io_rdAddr_2; // @[LVTMultiPortRams.scala 52:21 LVTMultiPortRams.scala 60:30]
  assign Memory_5_io_wrEna = io_wrEna_1; // @[LVTMultiPortRams.scala 52:21 LVTMultiPortRams.scala 57:29]
  assign Memory_5_io_wrData = io_wrData_1; // @[LVTMultiPortRams.scala 52:21 LVTMultiPortRams.scala 59:30]
  assign Memory_5_io_wrAddr = io_wrAddr_1; // @[LVTMultiPortRams.scala 52:21 LVTMultiPortRams.scala 58:30]
  assign Memory_6_clock = clock;
  assign Memory_6_io_rdAddr = io_rdAddr_0; // @[LVTMultiPortRams.scala 52:21 LVTMultiPortRams.scala 60:30]
  assign Memory_6_io_wrEna = io_wrEna_2; // @[LVTMultiPortRams.scala 52:21 LVTMultiPortRams.scala 57:29]
  assign Memory_6_io_wrData = io_wrData_2; // @[LVTMultiPortRams.scala 52:21 LVTMultiPortRams.scala 59:30]
  assign Memory_6_io_wrAddr = io_wrAddr_2; // @[LVTMultiPortRams.scala 52:21 LVTMultiPortRams.scala 58:30]
  assign Memory_7_clock = clock;
  assign Memory_7_io_rdAddr = io_rdAddr_1; // @[LVTMultiPortRams.scala 52:21 LVTMultiPortRams.scala 60:30]
  assign Memory_7_io_wrEna = io_wrEna_2; // @[LVTMultiPortRams.scala 52:21 LVTMultiPortRams.scala 57:29]
  assign Memory_7_io_wrData = io_wrData_2; // @[LVTMultiPortRams.scala 52:21 LVTMultiPortRams.scala 59:30]
  assign Memory_7_io_wrAddr = io_wrAddr_2; // @[LVTMultiPortRams.scala 52:21 LVTMultiPortRams.scala 58:30]
  assign Memory_8_clock = clock;
  assign Memory_8_io_rdAddr = io_rdAddr_2; // @[LVTMultiPortRams.scala 52:21 LVTMultiPortRams.scala 60:30]
  assign Memory_8_io_wrEna = io_wrEna_2; // @[LVTMultiPortRams.scala 52:21 LVTMultiPortRams.scala 57:29]
  assign Memory_8_io_wrData = io_wrData_2; // @[LVTMultiPortRams.scala 52:21 LVTMultiPortRams.scala 59:30]
  assign Memory_8_io_wrAddr = io_wrAddr_2; // @[LVTMultiPortRams.scala 52:21 LVTMultiPortRams.scala 58:30]
  assign lvt_clock = clock;
  assign lvt_reset = reset;
  assign lvt_io_wrAddr_0 = io_wrAddr_0; // @[LVTMultiPortRams.scala 65:22]
  assign lvt_io_wrAddr_1 = io_wrAddr_1; // @[LVTMultiPortRams.scala 65:22]
  assign lvt_io_wrAddr_2 = io_wrAddr_2; // @[LVTMultiPortRams.scala 65:22]
  assign lvt_io_wrEna_0 = io_wrEna_0; // @[LVTMultiPortRams.scala 64:21]
  assign lvt_io_wrEna_1 = io_wrEna_1; // @[LVTMultiPortRams.scala 64:21]
  assign lvt_io_wrEna_2 = io_wrEna_2; // @[LVTMultiPortRams.scala 64:21]
  assign lvt_io_rdAddr_0 = io_rdAddr_0; // @[LVTMultiPortRams.scala 68:22]
  assign lvt_io_rdAddr_1 = io_rdAddr_1; // @[LVTMultiPortRams.scala 68:22]
  assign lvt_io_rdAddr_2 = io_rdAddr_2; // @[LVTMultiPortRams.scala 68:22]

  integer addr_0 = 4'h5;
  integer data_0 = 8'h1f;
  integer addr_1 = 4'h6;
  integer data_1 = 8'h7;
  integer addr_2 = 4'h7;
  integer data_2 = 8'h9;
  // multi-port
  sequence ant0;
    (reset == 0) && (io_wrAddr_0 == addr_0) && (io_wrData_0 == data_0) && (io_wrEna_0 == 1'b1) &&
    (io_wrAddr_1 == addr_1) && (io_wrData_1 == data_1) && (io_wrEna_1 == 1'b1) &&
    (io_wrAddr_2 == addr_2) && (io_wrData_2 == data_2) && (io_wrEna_2 == 1'b1);
  endsequence
  sequence u0;
    ##1 (lvt.lvtReg_5 == 0) && (Memory.mem[5] == data_0) && (Memory_1.mem[5] == data_0) && (Memory_2.mem[5] == data_0) 
    && (lvt.lvtReg_6 == 1) && (Memory_3.mem[6] == data_1) && (Memory_4.mem[6] == data_1)&& (Memory_5.mem[6] == data_1)
    && (lvt.lvtReg_7 == 2) && (Memory_6.mem[7] == data_2) && (Memory_7.mem[7] == data_2)&& (Memory_8.mem[7] == data_2);
  endsequence
  assert property(@(posedge clock) ant0 |-> u0);

  sequence ant1;
    ((reset == 0) &&  (lvt.lvtReg_5 == 0) && (Memory.mem[5] == data_0) && (Memory_1.mem[5] == data_0) && (Memory_2.mem[5] == data_0) 
    && (lvt.lvtReg_6 == 1) && (Memory_3.mem[6] == data_1) && (Memory_4.mem[6] == data_1)&& (Memory_5.mem[6] == data_1)
    && (lvt.lvtReg_7 == 2) && (Memory_6.mem[7] == data_2) && (Memory_7.mem[7] == data_2)&& (Memory_8.mem[7] == data_2)
    && (io_wrEna_0 == 1'b0 || (io_wrAddr_0 != addr_0 && io_wrAddr_0 != addr_1 && io_wrAddr_0 != addr_2)) 
    && (io_wrEna_1 == 1'b0 || (io_wrAddr_1 != addr_0 && io_wrAddr_1 != addr_1 &&io_wrAddr_1 != addr_2))
    && (io_wrEna_2 == 1'b0 || (io_wrAddr_2 != addr_0 && io_wrAddr_2 != addr_1 &&io_wrAddr_2 != addr_2))) 
    ##1 ((reset == 0) && (io_wrEna_0 == 1'b0 || (io_wrAddr_0 != addr_0 && io_wrAddr_0 != addr_1 && io_wrAddr_0 != addr_2)) 
    && (io_wrEna_1 == 1'b0 || (io_wrAddr_1 != addr_0 && io_wrAddr_1 != addr_1 &&io_wrAddr_1 != addr_2))
    && (io_wrEna_2 == 1'b0 || (io_wrAddr_2 != addr_0 && io_wrAddr_2 != addr_1 &&io_wrAddr_2 != addr_2)))[*3];
  endsequence
  sequence u1;
    ##1 (lvt.lvtReg_5 == 0) && (Memory.mem[5] == data_0) && (Memory_1.mem[5] == data_0) && (Memory_2.mem[5] == data_0) 
    && (lvt.lvtReg_6 == 1) && (Memory_3.mem[6] == data_1) && (Memory_4.mem[6] == data_1)&& (Memory_5.mem[6] == data_1)
    && (lvt.lvtReg_7 == 2) && (Memory_6.mem[7] == data_2) && (Memory_7.mem[7] == data_2)&& (Memory_8.mem[7] == data_2);
  endsequence
  assert property(@(posedge clock) ant1 |-> u1);

  sequence ant2;
    (lvt.lvtReg_5 == 0) && (Memory.mem[5] == data_0) && (Memory_1.mem[5] == data_0) && (Memory_2.mem[5] == data_0) 
    && (lvt.lvtReg_6 == 1) && (Memory_3.mem[6] == data_1) && (Memory_4.mem[6] == data_1)&& (Memory_5.mem[6] == data_1)
    && (lvt.lvtReg_7 == 2) && (Memory_6.mem[7] == data_2) && (Memory_7.mem[7] == data_2)&& (Memory_8.mem[7] == data_2) &&
    (io_rdAddr_0 == addr_0) && (io_rdAddr_1 == addr_1) && (io_rdAddr_2 == addr_2) ;
  endsequence
  sequence cons2;
    (io_rdData_0 == data_0) && (io_rdData_1 == data_1) && (io_rdAddr_2 == addr_2);
  endsequence
  assert property(@(posedge clock) ant2 |-> cons2);
endmodule
